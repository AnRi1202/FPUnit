library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity FPMult_NoRA is
    port (clk : in std_logic;
          X : in  std_logic_vector(8+23+2 downto 0);
          Y : in  std_logic_vector(8+23+2 downto 0);
          R : out  std_logic_vector(8+23+2 downto 0);
         --  round_out : out std_logic;
         --  expSig_out : out std_logic_vector(32 downto 0);
         --  expSigPostRound_in : in std_logic_vector(32 downto 0);
          -- Shared IntAdder_27 ports for exp calculations
          expAdder_X_out : out std_logic_vector(7 downto 0);
          expAdder_Y_out : out std_logic_vector(7 downto 0);
          expAdder_Cin_out : out std_logic;
          expAdder_R_in : in std_logic_vector(26 downto 0) );
end entity;

architecture arch of FPMult_NoRA is 
   component IntMultiplier_24x24_48_Freq1_uid5 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(23 downto 0);
             Y : in  std_logic_vector(23 downto 0);
             R : out  std_logic_vector(47 downto 0)   );
   end component;

   component IntAdder_33_Freq1_uid280 is
      port ( clk : in std_logic;
             X : in  std_logic_vector(32 downto 0);
             Y : in  std_logic_vector(32 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(32 downto 0)   );
   end component;

signal sign :  std_logic;
   -- timing of sign: (c0, 0.043000ns)
signal expX :  std_logic_vector(7 downto 0);
   -- timing of expX: (c0, 0.000000ns)
signal expY :  std_logic_vector(7 downto 0);
   -- timing of expY: (c0, 0.000000ns)
signal expSumPreSub :  std_logic_vector(9 downto 0);
   -- timing of expSumPreSub: (c0, 1.092000ns)
signal bias :  std_logic_vector(9 downto 0);
   -- timing of bias: (c0, 0.000000ns)
signal expSum :  std_logic_vector(9 downto 0);
   -- timing of expSum: (c0, 2.184000ns)
signal sigX :  std_logic_vector(23 downto 0);
   -- timing of sigX: (c0, 0.000000ns)
signal sigY :  std_logic_vector(23 downto 0);
   -- timing of sigY: (c0, 0.000000ns)
signal sigProd :  std_logic_vector(47 downto 0);
   -- timing of sigProd: (c0, 4.870000ns)
   signal excSel :  std_logic_vector(3 downto 0);
   signal exc :  std_logic_vector(1 downto 0);
   signal norm :  std_logic;
   signal expPostNorm :  std_logic_vector(9 downto 0);
   signal sigProdExt :  std_logic_vector(47 downto 0);
   signal expSig :  std_logic_vector(32 downto 0);
   signal sticky :  std_logic;
   signal guard :  std_logic;
   signal round :  std_logic;
   signal expSigPostRound :  std_logic_vector(32 downto 0);
   signal excPostNorm :  std_logic_vector(1 downto 0);
   signal finalExc :  std_logic_vector(1 downto 0);
begin
   sign <= X(31) xor Y(31);
   expX <= X(30 downto 23);
   expY <= Y(30 downto 23);
   
   -- Use shared IntAdder_27 for expSumPreSub calculation
   -- Pad 10-bit values to 27-bit
   expAdder_X_out <=expX;  -- 8bit  
   expAdder_Y_out <=expY;  -- 8bit
   expAdder_Cin_out <= '0';
   expSumPreSub <= '0' & expAdder_R_in(8 downto 0);  -- Extract lower 10 bits
   
   bias <= CONV_STD_LOGIC_VECTOR(127,10);
   expSum <= expSumPreSub - bias;
   sigX <= "1" & X(22 downto 0);
   sigY <= "1" & Y(22 downto 0);
   SignificandMultiplication: IntMultiplier_24x24_48_Freq1_uid5
      port map ( clk  => clk,
                 X => sigX,
                 Y => sigY,
                 R => sigProd); -- 48bit
   excSel <= X(33 downto 32) & Y(33 downto 32);
   with excSel  select  
   exc <= "00" when  "0000" | "0001" | "0100", 
          "01" when "0101",
          "10" when "0110" | "1001" | "1010" ,
          "11" when others;

   norm <= sigProd(47); -- 最大桁
   -- exponent update
   expPostNorm <= expSum + ("000000000" & norm); -- 最上位が1ならexpを1つ挙げる. [1,2)同士の掛け算は[2,4), 11ならnormが1になるからexpを上げる
   -- significand normalization shift
   sigProdExt <= sigProd(46 downto 0) & "0" when norm='1' else
                         sigProd(45 downto 0) & "00"; --normが0なら01. . ってつづくから1でカットしていい
   expSig <= expPostNorm & sigProdExt(47 downto 25);
   sticky <= sigProdExt(24); -- addとは意味が違う sticky, guardの順番(addはguard, stickyだった)
   guard <= '0' when sigProdExt(23 downto 0)="000000000000000000000000" else '1';
   round <= sticky and ( (guard and not(sigProdExt(25))) or (sigProdExt(25) ))  ;
   RoundingAdder: IntAdder_33_Freq1_uid280
      port map ( clk  => clk,
                 Cin => round,
                 X => expSig,
                 Y => "000000000000000000000000000000000",
                 R => expSigPostRound);
   -- round_out <= round;
   -- expSig_out <= expSig;
   -- expSigPostRound <= expSigPostRound_in;

   with expSigPostRound(32 downto 31)  select 
   excPostNorm <=  "01"  when  "00",
                               "10"             when "01", 
                               "00"             when "11"|"10",
                               "11"             when others;
   with exc  select  
   finalExc <= exc when  "11"|"10"|"00",
                       excPostNorm when others; 
   R <= finalExc & sign & expSigPostRound(30 downto 0);
end architecture;
