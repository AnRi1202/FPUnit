library ieee;
use ieee.std_logic_1164.all;

entity tb_fpsqrt_kintex is
end tb_fpsqrt_kintex;



