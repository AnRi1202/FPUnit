../src_shared_combine_sv/FPALL_pkg.sv