module tb_FPALL_shared;


endmodule